module stage_MEM ();



endmodule
