module EX_stage();


  
endmodule
