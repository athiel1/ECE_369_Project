module stage_ID ();



endmodule
