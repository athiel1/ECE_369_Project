module stage_EX ();



endmodule
