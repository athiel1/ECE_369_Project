module stage_IF ();
    input 


endmodule
