module stage_WB ();



endmodule
