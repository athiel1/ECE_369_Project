module stage_IF ();



endmodule
